// Name : Gaurang Pandey
// File : snn_core.sv
// Description : 
//


module snn_core;

  // This is a placeholder file

endmodule 
