// Name : Gaurang Pandey
// File : top.sv
// Description :
//


module top;

  // This is placeholder

endmodule
