// List of the SNN sequences

`include "snn_base_sequence.sv"
`include "snn_reg_rand_sequence.sv"
`include "snn_reg_bitbash_sequence.sv"
`include "snn_init_sequence.sv"
`include "snn_stripe_sequence.sv"
`include "snn_digit_sequence.sv"
`include "snn_checkered_sequence.sv"
`include "snn_gradient_sequence.sv"
`include "snn_radial_sequence.sv"
`include "snn_noise_pattern_sequence.sv"
`include "snn_random_sequence.sv"