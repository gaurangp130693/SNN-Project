// List of the SNN sequences

`include "snn_base_sequence.sv"
`include "snn_init_sequence.sv"
`include "snn_pixel_sequence.sv"